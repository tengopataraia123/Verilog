module alu(
	input [31:0] A_in,
	input [31:0] B_in,
	input [3:0] cmd_in,
	input [1:0] sh_in,
	input [4:0] shamt5_in,
	input I_in,
	input S_in,

	output [31:0] Result_out,
	output [3:0] NZCV_out);
	
	reg [32:0] result = 0;
	reg [3:0] NZCV = 0;
	
	assign Result_out[31:0] = result[31:0];
	assign NZCV_out = NZCV;
	
	always@(*) begin
		
	end
	
endmodule 